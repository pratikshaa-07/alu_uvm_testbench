package pkg;
  import uvm_pkg::*;
`include "uvm_macros.svh"
`include "item.sv"
`include "seq.sv"
`include "seqr.sv"
`include "drv.sv"
`include "mon.sv"
`include "agt.sv"
`include "sb.sv"
`include "cov.sv"
`include "env.sv"
`include "test.sv"
endpackage
