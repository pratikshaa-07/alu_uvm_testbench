package pkg;
`include "uvm_pkg.sv"
`include "uvm_macros.svh"
`include "item.sv"
`include "seq.sv"
`include "seqr.sv"
`include "drv.sv"
`include "mon.sv"
`include "agt.sv"
`include "sb.sv"
`include "covg.sv"
`include "env.sv"
`include "tb.sv"
endpackage
