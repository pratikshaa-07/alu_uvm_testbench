`define oplen 8
`define cmdlen 4
